//-----------------------------------------------------------------------------
// Company    : u-blox Cork, Ireland
// Created    : Monday, 02 March 2015 08:48PM
// Last commit: $Date: 2015/06/04 $
// Updated by : $Author: prya $
//-----------------------------------------------------------------------------
// Copyright (c) 2014 u-blox Cork, Ireland
//-----------------------------------------------------------------------------
// $Id: //depot/icm/proj/ic_mx_dig_top/trunk/rtl/mx_dig_top/mx_apb_mmap.v#5 $
// AUTO-GENERATED: Do Not Hand Edit
//-----------------------------------------------------------------------------

module mx_apb_mmap(
  input sig1,sig2, sig3,            // these types of ports don't work yet
  sig4, sig5;
	input   wire                PClkxCI,
	input                   PResetxARBI,
	output reg              PEnClkxSO,
	input                   PEnClkxSI,
	input           [31:0]  PAddrxDI,
	input                   PSelxSI,
	input                   PEnablexSI,
	input                   PWritexSI,
	input           [31:0]  PWDataxDI,
	output  reg             PReadyxSO,
	output  reg     [31:0]  PRDataxDO,
	output  reg             PSlverrxSO,
	output                  Meas_ldoBypassxO,           // this is a comment
	output                  Meas_ldoEnablexO,/// I'm a comment too
// I'm just in the way  
	output                  Meas_ldoFast_lockxO,
	input           [15:0]  Hist_q_5Hist_out_i_10xI,
	input /*important shit to be said*/          [15:0]  Hist_q_5Hist_out_i_11xI,
	input           [15:0]  Hist_q_6Hist_out_i_12xI,
	input           [15:0]  Hist_q_6Hist_out_i_13xI,
  /* howa
   * about 
   here then
   adsf */
	input           [15:0]  Hist_q_7Hist_out_i_14xI,
	input           [15:0]  Hist_q_7Hist_out_i_15xI,
	input           [15:0]  Hist_q_8Hist_out_i_16xI,
	input           [15:0]  Hist_q_8Hist_out_i_17xI,
	input           [15:0]  Hist_q_9Hist_out_i_18xI,
/*asdf*/

	input           [15:0]  Hist_q_9Hist_out_i_19xI,
	input           [15:0]  Hist_q_10Hist_out_i_20xI,
	input           [15:0]  Hist_q_10Hist_out_i_21xI,
	input           [15:0]  Hist_q_11Hist_out_i_22xI,input           [15:0]  Hist_q_11Hist_out_i_23xI,
	input           [15:0]  Hist_q_12Hist_out_i_24xI,	input           [15:0]  Hist_q_12Hist_out_i_25xI,
	input           [15:0]  Hist_q_13Hist_out_i_26xI,
	input           [15:0]  Hist_q_13Hist_out_i_27xI,
	input           [15:0]  Hist_q_14Hist_out_i_28xI,
	input           [15:0]  Hist_q_14Hist_out_i_29xI,
	input           [15:0]  Hist_q_15Hist_out_i_30xI,
	input           [15:0]  Hist_q_15Hist_out_i_31xI,output           [3:0]  Adc_tmodeTmodexO
  );

  reg           PSelxSI_meas;
  reg           PSelxSI_measADC;
  reg           PSelxSI_measADCflags;
  reg           PSelxSI_measDFE;
 
  wire          PEnClkxSO_meas, PEnClkxSO_measADC, PEnClkxSO_measDFE, PEnClkxSO_measADCflags;
  wire          PReadyxSO_meas, PReadyxSO_measADC, PReadyxSO_measDFE, PReadyxSO_measADCflags;
  wire [31:0]   PRDataxDO_meas, PRDataxDO_measADC, PRDataxDO_measDFE, PRDataxDO_measADCflags;
  wire          PSlverrxSO_meas, PSlverrxSO_measADC, PSlverrxSO_measDFE, PSlverrxSO_measADCflags;

// Sel decode for the each block
always @*
  begin

  PSelxSI_meas         = 1'b0;
  PSelxSI_measADC      = 1'b0;
  PSelxSI_measADCflags = 1'b0;
  PSelxSI_measDFE      = 1'b0;
  PEnClkxSO            = 1'b0;
  PReadyxSO            = 1'b0;
  PRDataxDO            = 32'h0;
  PSlverrxSO           = 1'b0;

  if(PSelxSI) begin
    PEnClkxSO  = PEnClkxSO_meas | PEnClkxSO_measADC | PEnClkxSO_measDFE | PEnClkxSO_measADCflags;
    PReadyxSO  = PReadyxSO_meas & PReadyxSO_measADC & PReadyxSO_measDFE & PReadyxSO_measADCflags;
    PSlverrxSO = PSlverrxSO_meas| PSlverrxSO_measADC| PSlverrxSO_measDFE| PSlverrxSO_measADCflags;
  end 

  case(PAddrxDI[12:11])
    2'b00:  begin
      PSelxSI_meas         = PSelxSI;
      PRDataxDO            = PRDataxDO_meas;
    end
    2'b01:  begin
      PSelxSI_measADC      = PSelxSI;
      PRDataxDO            = PRDataxDO_measADC;
    end
    2'b10:  begin
      PSelxSI_measDFE      = PSelxSI;
      PRDataxDO            = PRDataxDO_measDFE;
    end
    2'b11:  begin  
      PSelxSI_measADCflags = PSelxSI;
      PRDataxDO            = PRDataxDO_measADCflags;
    end
  endcase
  end

mx_apb_mmap_meas mx_apb_mmap_meas (
    .PClkxCI                                   (PClkxCI),
    .PResetxARBI                               (PResetxARBI),
    .PEnClkxSO                                 (PEnClkxSO_meas),
    .PEnClkxSI                                 (PEnClkxSI),
    .PAddrxDI                                  ({21'h0, PAddrxDI[10:0]}),
    .PSelxSI                                   (PSelxSI_meas),
    .PEnablexSI                                (PEnablexSI),
    .PWritexSI                                 (PWritexSI),
    .PWDataxDI                                 (PWDataxDI),
    .PReadyxSO                                 (PReadyxSO_meas),
    .PRDataxDO                                 (PRDataxDO_meas),
    .PSlverrxSO                                (PSlverrxSO_meas),
    .Meas_ldoBypassxO                          (Meas_ldoBypassxO),
    .Meas_ldoEnablexO                          (Meas_ldoEnablexO),
    .Meas_ldoFast_lockxO                       (Meas_ldoFast_lockxO),
    .Meas_ldoVout_ctrlxO                       (Meas_ldoVout_ctrlxO),
    .Adc_ldoBypassxO                           (Adc_ldoBypassxO),
    .Adc_ldoEnablexO                           (Adc_ldoEnablexO),
    .Adc_ldoFast_lockxO                        (Adc_ldoFast_lockxO),
    .Adc_ldoVout_ctrlxO                        (Adc_ldoVout_ctrlxO),
    .Cal_ldoBypassxO                           (Cal_ldoBypassxO),
    .Cal_ldoEnablexO                           (Cal_ldoEnablexO),
    .Cal_ldoFast_lockxO                        (Cal_ldoFast_lockxO),
    .Cal_ldoVout_ctrlxO                        (Cal_ldoVout_ctrlxO),
    .MeasRxrf_enxO                             (MeasRxrf_enxO),
    .MeasSf_enxO                               (MeasSf_enxO),
    .MeasDac_enxO                              (MeasDac_enxO),
    .MeasDiv_enxO                              (MeasDiv_enxO),
    .MeasTempcell_enxO                         (MeasTempcell_enxO),
    .MeasMeas_cal_enxO                         (MeasMeas_cal_enxO),
    .MeasBypxO                                 (MeasBypxO),
    .MeasSelxO                                 (MeasSelxO),
    .MeasIqmuxxO                               (MeasIqmuxxO),
    .MeasClkgen_enxO                           (MeasClkgen_enxO),
    .EnablesAdc_i_enxO                         (EnablesAdc_i_enxO),
    .EnablesAdc_q_enxO                         (EnablesAdc_q_enxO),
    .Meas_gainGtrimxO                          (Meas_gainGtrimxO),
    .Meas_gainLna_rxO                          (Meas_gainLna_rxO),
    .Meas_gainAttxO                            (Meas_gainAttxO),
    .Meas_tfCtrimxO                            (Meas_tfCtrimxO),
    .Meas_dacPixO                              (Meas_dacPixO),
    .Meas_dacNixO                              (Meas_dacNixO),
    .Meas_dacPqxO                              (Meas_dacPqxO),
    .Meas_dacNqxO                              (Meas_dacNqxO),
    .ClkgenMod_pxO                             (ClkgenMod_pxO),
    .CalEnxO                                   (CalEnxO),
    .CalIbiasxO                                (CalIbiasxO),
    .CalConstgmxO                              (CalConstgmxO),
    .Cal_gainGmxO                              (Cal_gainGmxO),
    .Cal_gainFbxO                              (Cal_gainFbxO),
    .Cal_gainCasnxO                            (Cal_gainCasnxO),
    .Cal_gainCaspxO                            (Cal_gainCaspxO),
    .AtstMeas_en_AxO                           (AtstMeas_en_AxO),
    .AtstMeas_en_BxO                           (AtstMeas_en_BxO),
    .AtstMeas_en_CxO                           (AtstMeas_en_CxO),
    .AtstMeas_en_DxO                           (AtstMeas_en_DxO),
    .AtstMeas_en_ExO                           (AtstMeas_en_ExO),
    .AtstMeas_en_FxO                           (AtstMeas_en_FxO),
    .AtstMeas_ldo_en_AxO                       (AtstMeas_ldo_en_AxO),
    .AtstAdc_ldo_en_AxO                        (AtstAdc_ldo_en_AxO),
    .AtstCal_en_AxO                            (AtstCal_en_AxO),
    .AtstCal_en_BxO                            (AtstCal_en_BxO),
    .AtstCal_en_CxO                            (AtstCal_en_CxO),
    .AtstCal_ldo_en_AxO                        (AtstCal_ldo_en_AxO),
    .AtstAdc_i_en_AxO                          (AtstAdc_i_en_AxO),
    .AtstAdc_i_en_BxO                          (AtstAdc_i_en_BxO),
    .AtstAdc_q_en_AxO                          (AtstAdc_q_en_AxO),
    .AtstAdc_q_en_BxO                          (AtstAdc_q_en_BxO),
    .Atst_toplevelMeas_en_AxO                  (Atst_toplevelMeas_en_AxO),
    .Atst_toplevelMeas_en_BxO                  (Atst_toplevelMeas_en_BxO),
    .Atst_toplevelMeas_en_CxO                  (Atst_toplevelMeas_en_CxO),
    .Atst_toplevelMeas_en_DxO                  (Atst_toplevelMeas_en_DxO),
    .Atst_toplevelMeas_en_ExO                  (Atst_toplevelMeas_en_ExO),
    .Atst_toplevelMeas_en_FxO                  (Atst_toplevelMeas_en_FxO),
    .Atst_toplevelMeas_ldo_en_AxO              (Atst_toplevelMeas_ldo_en_AxO),
    .Atst_toplevelAdc_ldo_en_AxO               (Atst_toplevelAdc_ldo_en_AxO),
    .Atst_toplevelCal_en_AxO                   (Atst_toplevelCal_en_AxO),
    .Atst_toplevelCal_en_BxO                   (Atst_toplevelCal_en_BxO),
    .Atst_toplevelCal_en_CxO                   (Atst_toplevelCal_en_CxO),
    .Atst_toplevelCal_ldo_en_AxO               (Atst_toplevelCal_ldo_en_AxO),
    .Atst_toplevelAdc_i_en_AxO                 (Atst_toplevelAdc_i_en_AxO),
    .Atst_toplevelAdc_i_en_BxO                 (Atst_toplevelAdc_i_en_BxO),
    .Atst_toplevelAdc_q_en_AxO                 (Atst_toplevelAdc_q_en_AxO),
    .Atst_toplevelAdc_q_en_BxO                 (Atst_toplevelAdc_q_en_BxO),
    .Adc_clkMuxClkin_selxO                     (Adc_clkMuxClkin_selxO),
    .Adc_clkMuxAdc_clk_selxO                   (Adc_clkMuxAdc_clk_selxO),
    .Adc_clkMuxDig_clk_selxO                   (Adc_clkMuxDig_clk_selxO),
    .Adc_clkMuxTx_clk_selxO                    (Adc_clkMuxTx_clk_selxO),
    .Adc_clkMuxAdc_dfe_clk_invertxO            (Adc_clkMuxAdc_dfe_clk_invertxO),
    .Meas_spareMainxO                          (Meas_spareMainxO),
    .Meas_spareIxO                             (Meas_spareIxO),
    .Meas_spareQxO                             (Meas_spareQxO),
    .Cal_spareMainxO                           (Cal_spareMainxO),
    .Atst_measMaster_enxO                      (Atst_measMaster_enxO),
    .Atst_measMaster_pulldownxO                (Atst_measMaster_pulldownxO),
    .Atst_measAuxAdc_enxO                      (Atst_measAuxAdc_enxO)
  );

mx_apb_mmap_measADC mx_apb_mmap_measADC (
    .PClkxCI                                   (PClkxCI),
    .PResetxARBI                               (PResetxARBI),
    .PEnClkxSO                                 (PEnClkxSO_measADC),
    .PEnClkxSI                                 (PEnClkxSI),
    .PAddrxDI                                  ({21'h0, PAddrxDI[10:0]}),
    .PSelxSI                                   (PSelxSI_measADC),
    .PEnablexSI                                (PEnablexSI),
    .PWritexSI                                 (PWritexSI),
    .PWDataxDI                                 (PWDataxDI),
    .PReadyxSO                                 (PReadyxSO_measADC),
    .PRDataxDO                                 (PRDataxDO_measADC),
    .PSlverrxSO                                (PSlverrxSO_measADC),
    .Adc_mode_iAdcModexO                       (Adc_mode_iAdcModexO),
    .Adc_mode_iInterleaveModexO                (Adc_mode_iInterleaveModexO),
    .Adc_mode_iCH1enxO                         (Adc_mode_iCH1enxO),
    .Adc_mode_iCH2enxO                         (Adc_mode_iCH2enxO),
    .Adc_mode_qAdcModexO                       (Adc_mode_qAdcModexO),
    .Adc_mode_qInterleaveModexO                (Adc_mode_qInterleaveModexO),
    .Adc_mode_qCH1enxO                         (Adc_mode_qCH1enxO),
    .Adc_mode_qCH2enxO                         (Adc_mode_qCH2enxO),
    .Adc_cal_statusCHI1OfflineCalDonexI        (Adc_cal_statusCHI1OfflineCalDonexI),
    .Adc_cal_statusCHI2OfflineCalDonexI        (Adc_cal_statusCHI2OfflineCalDonexI),
    .Adc_cal_statusCHQ1OfflineCalDonexI        (Adc_cal_statusCHQ1OfflineCalDonexI),
    .Adc_cal_statusCHQ2OfflineCalDonexI        (Adc_cal_statusCHQ2OfflineCalDonexI),
    .Adc_i_calclkCalClkDivxO                   (Adc_i_calclkCalClkDivxO),
    .Adc_q_calclkCalClkDivxO                   (Adc_q_calclkCalClkDivxO),
    .Adc_i_ditherDitherEnxO                    (Adc_i_ditherDitherEnxO),
    .Adc_i_ditherDitherRevertxO                (Adc_i_ditherDitherRevertxO),
    .Adc_i_ditherDitherDelayxO                 (Adc_i_ditherDitherDelayxO),
    .Adc_q_ditherDitherEnxO                    (Adc_q_ditherDitherEnxO),
    .Adc_q_ditherDitherRevertxO                (Adc_q_ditherDitherRevertxO),
    .Adc_q_ditherDitherDelayxO                 (Adc_q_ditherDitherDelayxO),
    .Adc_iqmuxEn_ixO                           (Adc_iqmuxEn_ixO),
    .Adc_iqmuxEn_qxO                           (Adc_iqmuxEn_qxO),
    .Adc_cal_readback_ctrlSelectIxO            (Adc_cal_readback_ctrlSelectIxO),
    .Adc_cal_readback_ctrlSelectQxO            (Adc_cal_readback_ctrlSelectQxO),
    .Adc_cal_readback_iResultxI                (Adc_cal_readback_iResultxI),
    .Adc_cal_readback_qResultxI                (Adc_cal_readback_qResultxI),
    .CHI1_calCH1calModexO                      (CHI1_calCH1calModexO),
    .CHI1_calShortADCInputxO                   (CHI1_calShortADCInputxO),
    .CHI1_calStageCtrlStageDisablexO           (CHI1_calStageCtrlStageDisablexO),
    .CHI1_ChannelGainCH1channelGainxO          (CHI1_ChannelGainCH1channelGainxO),
    .CHI1_DACN1CH1capControlN1xO               (CHI1_DACN1CH1capControlN1xO),
    .CHI1_DACP1CH1capControlP1xO               (CHI1_DACP1CH1capControlP1xO),
    .CHI1_DACN2CH1capControlN2xO               (CHI1_DACN2CH1capControlN2xO),
    .CHI1_DACP2CH1capControlP2xO               (CHI1_DACP2CH1capControlP2xO),
    .CHI1_AMPCH1AmpGainCalPxO                  (CHI1_AMPCH1AmpGainCalPxO),
    .CHI1_AMPCH1AmpGainCalNxO                  (CHI1_AMPCH1AmpGainCalNxO),
    .CHI1_AMPCH1increaseAmpDelayxO             (CHI1_AMPCH1increaseAmpDelayxO),
    .CHI1_MSBCALCH1MSBCalxO                    (CHI1_MSBCALCH1MSBCalxO),
    .CHI1_comp12CalPComp_calxO                 (CHI1_comp12CalPComp_calxO),
    .CHI1_comp12CalNComp_calxO                 (CHI1_comp12CalNComp_calxO),
    .CHI1_comp11CalPComp_calxO                 (CHI1_comp11CalPComp_calxO),
    .CHI1_comp11CalNComp_calxO                 (CHI1_comp11CalNComp_calxO),
    .CHI1_comp10CalPComp_calxO                 (CHI1_comp10CalPComp_calxO),
    .CHI1_comp10CalNComp_calxO                 (CHI1_comp10CalNComp_calxO),
    .CHI1_comp9CalPComp_calxO                  (CHI1_comp9CalPComp_calxO),
    .CHI1_comp9CalNComp_calxO                  (CHI1_comp9CalNComp_calxO),
    .CHI1_comp8CalPComp_calxO                  (CHI1_comp8CalPComp_calxO),
    .CHI1_comp8CalNComp_calxO                  (CHI1_comp8CalNComp_calxO),
    .CHI1_comp7CalPComp_calxO                  (CHI1_comp7CalPComp_calxO),
    .CHI1_comp7CalNComp_calxO                  (CHI1_comp7CalNComp_calxO),
    .CHI1_comp6CalPComp_calxO                  (CHI1_comp6CalPComp_calxO),
    .CHI1_comp6CalNComp_calxO                  (CHI1_comp6CalNComp_calxO),
    .CHI1_comp5CalPComp_calxO                  (CHI1_comp5CalPComp_calxO),
    .CHI1_comp5CalNComp_calxO                  (CHI1_comp5CalNComp_calxO),
    .CHI1_comp4CalPComp_calxO                  (CHI1_comp4CalPComp_calxO),
    .CHI1_comp4CalNComp_calxO                  (CHI1_comp4CalNComp_calxO),
    .CHI1_comp3CalPComp_calxO                  (CHI1_comp3CalPComp_calxO),
    .CHI1_comp3CalNComp_calxO                  (CHI1_comp3CalNComp_calxO),
    .CHI1_comp2CalPComp_calxO                  (CHI1_comp2CalPComp_calxO),
    .CHI1_comp2CalNComp_calxO                  (CHI1_comp2CalNComp_calxO),
    .CHI1_comp1CalPComp_calxO                  (CHI1_comp1CalPComp_calxO),
    .CHI1_comp1CalNComp_calxO                  (CHI1_comp1CalNComp_calxO),
    .CHI1_comp0CalPComp_calxO                  (CHI1_comp0CalPComp_calxO),
    .CHI1_comp0CalNComp_calxO                  (CHI1_comp0CalNComp_calxO),
    .CHI1_compDelayCompDelayxO                 (CHI1_compDelayCompDelayxO),
    .CHI1_Fail_detectCH1p1CompFailFlagxI       (CHI1_Fail_detectCH1p1CompFailFlagxI),
    .CHI1_Fail_detectCH1p2CompFailFlagxI       (CHI1_Fail_detectCH1p2CompFailFlagxI),
    .CHI1_Fail_detectCH1AmpFailFlagxI          (CHI1_Fail_detectCH1AmpFailFlagxI),
    .CHI1_SPARESparexO                         (CHI1_SPARESparexO),
    .CHI1_N_ValuesNxO                          (CHI1_N_ValuesNxO),
    .CHI1_N_ValuesN2xO                         (CHI1_N_ValuesN2xO),
    .CHI1_N_ValuesN4xO                         (CHI1_N_ValuesN4xO),
    .CHI1_threshold12ThresholdxO               (CHI1_threshold12ThresholdxO),
    .CHI1_threshold11ThresholdxO               (CHI1_threshold11ThresholdxO),
    .CHI1_threshold10ThresholdxO               (CHI1_threshold10ThresholdxO),
    .CHI1_threshold9ThresholdxO                (CHI1_threshold9ThresholdxO),
    .CHI1_threshold8ThresholdxO                (CHI1_threshold8ThresholdxO),
    .CHI1_threshold7ThresholdxO                (CHI1_threshold7ThresholdxO),
    .CHI1_threshold6ThresholdxO                (CHI1_threshold6ThresholdxO),
    .CHI1_threshold5ThresholdxO                (CHI1_threshold5ThresholdxO),
    .CHI1_threshold4ThresholdxO                (CHI1_threshold4ThresholdxO),
    .CHI1_threshold3ThresholdxO                (CHI1_threshold3ThresholdxO),
    .CHI1_threshold2ThresholdxO                (CHI1_threshold2ThresholdxO),
    .CHI2_calCH2calModexO                      (CHI2_calCH2calModexO),
    .CHI2_calShortADCInputxO                   (CHI2_calShortADCInputxO),
    .CHI2_calStageCtrlStageDisablexO           (CHI2_calStageCtrlStageDisablexO),
    .CHI2_ChannelGainCH2channelGainxO          (CHI2_ChannelGainCH2channelGainxO),
    .CHI2_DACN1CH2capControlN1xO               (CHI2_DACN1CH2capControlN1xO),
    .CHI2_DACP1CH2capControlP1xO               (CHI2_DACP1CH2capControlP1xO),
    .CHI2_DACN2CH2capControlN2xO               (CHI2_DACN2CH2capControlN2xO),
    .CHI2_DACP2CH2capControlP2xO               (CHI2_DACP2CH2capControlP2xO),
    .CHI2_AMPCH2AmpGainCalPxO                  (CHI2_AMPCH2AmpGainCalPxO),
    .CHI2_AMPCH2AmpGainCalNxO                  (CHI2_AMPCH2AmpGainCalNxO),
    .CHI2_AMPCH2increaseAmpDelayxO             (CHI2_AMPCH2increaseAmpDelayxO),
    .CHI2_MSBCALCH2MSBCalxO                    (CHI2_MSBCALCH2MSBCalxO),
    .CHI2_comp12CalPComp_calxO                 (CHI2_comp12CalPComp_calxO),
    .CHI2_comp12CalNComp_calxO                 (CHI2_comp12CalNComp_calxO),
    .CHI2_comp11CalPComp_calxO                 (CHI2_comp11CalPComp_calxO),
    .CHI2_comp11CalNComp_calxO                 (CHI2_comp11CalNComp_calxO),
    .CHI2_comp10CalPComp_calxO                 (CHI2_comp10CalPComp_calxO),
    .CHI2_comp10CalNComp_calxO                 (CHI2_comp10CalNComp_calxO),
    .CHI2_comp9CalPComp_calxO                  (CHI2_comp9CalPComp_calxO),
    .CHI2_comp9CalNComp_calxO                  (CHI2_comp9CalNComp_calxO),
    .CHI2_comp8CalPComp_calxO                  (CHI2_comp8CalPComp_calxO),
    .CHI2_comp8CalNComp_calxO                  (CHI2_comp8CalNComp_calxO),
    .CHI2_comp7CalPComp_calxO                  (CHI2_comp7CalPComp_calxO),
    .CHI2_comp7CalNComp_calxO                  (CHI2_comp7CalNComp_calxO),
    .CHI2_comp6CalPComp_calxO                  (CHI2_comp6CalPComp_calxO),
    .CHI2_comp6CalNComp_calxO                  (CHI2_comp6CalNComp_calxO),
    .CHI2_comp5CalPComp_calxO                  (CHI2_comp5CalPComp_calxO),
    .CHI2_comp5CalNComp_calxO                  (CHI2_comp5CalNComp_calxO),
    .CHI2_comp4CalPComp_calxO                  (CHI2_comp4CalPComp_calxO),
    .CHI2_comp4CalNComp_calxO                  (CHI2_comp4CalNComp_calxO),
    .CHI2_comp3CalPComp_calxO                  (CHI2_comp3CalPComp_calxO),
    .CHI2_comp3CalNComp_calxO                  (CHI2_comp3CalNComp_calxO),
    .CHI2_comp2CalPComp_calxO                  (CHI2_comp2CalPComp_calxO),
    .CHI2_comp2CalNComp_calxO                  (CHI2_comp2CalNComp_calxO),
    .CHI2_comp1CalPComp_calxO                  (CHI2_comp1CalPComp_calxO),
    .CHI2_comp1CalNComp_calxO                  (CHI2_comp1CalNComp_calxO),
    .CHI2_comp0CalPComp_calxO                  (CHI2_comp0CalPComp_calxO),
    .CHI2_comp0CalNComp_calxO                  (CHI2_comp0CalNComp_calxO),
    .CHI2_compDelayCompDelayxO                 (CHI2_compDelayCompDelayxO),
    .CHI2_Fail_detectCH2p1CompFailFlagxI       (CHI2_Fail_detectCH2p1CompFailFlagxI),
    .CHI2_Fail_detectCH2p2CompFailFlagxI       (CHI2_Fail_detectCH2p2CompFailFlagxI),
    .CHI2_Fail_detectCH2AmpFailFlagxI          (CHI2_Fail_detectCH2AmpFailFlagxI),
    .CHI2_SPARESparexO                         (CHI2_SPARESparexO),
    .CHI2_N_ValuesNxO                          (CHI2_N_ValuesNxO),
    .CHI2_N_ValuesN2xO                         (CHI2_N_ValuesN2xO),
    .CHI2_N_ValuesN4xO                         (CHI2_N_ValuesN4xO),
    .CHI2_threshold12ThresholdxO               (CHI2_threshold12ThresholdxO),
    .CHI2_threshold11ThresholdxO               (CHI2_threshold11ThresholdxO),
    .CHI2_threshold10ThresholdxO               (CHI2_threshold10ThresholdxO),
    .CHI2_threshold9ThresholdxO                (CHI2_threshold9ThresholdxO),
    .CHI2_threshold8ThresholdxO                (CHI2_threshold8ThresholdxO),
    .CHI2_threshold7ThresholdxO                (CHI2_threshold7ThresholdxO),
    .CHI2_threshold6ThresholdxO                (CHI2_threshold6ThresholdxO),
    .CHI2_threshold5ThresholdxO                (CHI2_threshold5ThresholdxO),
    .CHI2_threshold4ThresholdxO                (CHI2_threshold4ThresholdxO),
    .CHI2_threshold3ThresholdxO                (CHI2_threshold3ThresholdxO),
    .CHI2_threshold2ThresholdxO                (CHI2_threshold2ThresholdxO),
    .CHQ1_calCH1calModexO                      (CHQ1_calCH1calModexO),
    .CHQ1_calShortADCInputxO                   (CHQ1_calShortADCInputxO),
    .CHQ1_calStageCtrlStageDisablexO           (CHQ1_calStageCtrlStageDisablexO),
    .CHQ1_ChannelGainCH1channelGainxO          (CHQ1_ChannelGainCH1channelGainxO),
    .CHQ1_DACN1CH1capControlN1xO               (CHQ1_DACN1CH1capControlN1xO),
    .CHQ1_DACP1CH1capControlP1xO               (CHQ1_DACP1CH1capControlP1xO),
    .CHQ1_DACN2CH1capControlN2xO               (CHQ1_DACN2CH1capControlN2xO),
    .CHQ1_DACP2CH1capControlP2xO               (CHQ1_DACP2CH1capControlP2xO),
    .CHQ1_AMPCH1AmpGainCalPxO                  (CHQ1_AMPCH1AmpGainCalPxO),
    .CHQ1_AMPCH1AmpGainCalNxO                  (CHQ1_AMPCH1AmpGainCalNxO),
    .CHQ1_AMPCH1increaseAmpDelayxO             (CHQ1_AMPCH1increaseAmpDelayxO),
    .CHQ1_MSBCALCH1MSBCalxO                    (CHQ1_MSBCALCH1MSBCalxO),
    .CHQ1_comp12CalPComp_calxO                 (CHQ1_comp12CalPComp_calxO),
    .CHQ1_comp12CalNComp_calxO                 (CHQ1_comp12CalNComp_calxO),
    .CHQ1_comp11CalPComp_calxO                 (CHQ1_comp11CalPComp_calxO),
    .CHQ1_comp11CalNComp_calxO                 (CHQ1_comp11CalNComp_calxO),
    .CHQ1_comp10CalPComp_calxO                 (CHQ1_comp10CalPComp_calxO),
    .CHQ1_comp10CalNComp_calxO                 (CHQ1_comp10CalNComp_calxO),
    .CHQ1_comp9CalPComp_calxO                  (CHQ1_comp9CalPComp_calxO),
    .CHQ1_comp9CalNComp_calxO                  (CHQ1_comp9CalNComp_calxO),
    .CHQ1_comp8CalPComp_calxO                  (CHQ1_comp8CalPComp_calxO),
    .CHQ1_comp8CalNComp_calxO                  (CHQ1_comp8CalNComp_calxO),
    .CHQ1_comp7CalPComp_calxO                  (CHQ1_comp7CalPComp_calxO),
    .CHQ1_comp7CalNComp_calxO                  (CHQ1_comp7CalNComp_calxO),
    .CHQ1_comp6CalPComp_calxO                  (CHQ1_comp6CalPComp_calxO),
    .CHQ1_comp6CalNComp_calxO                  (CHQ1_comp6CalNComp_calxO),
    .CHQ1_comp5CalPComp_calxO                  (CHQ1_comp5CalPComp_calxO),
    .CHQ1_comp5CalNComp_calxO                  (CHQ1_comp5CalNComp_calxO),
    .CHQ1_comp4CalPComp_calxO                  (CHQ1_comp4CalPComp_calxO),
    .CHQ1_comp4CalNComp_calxO                  (CHQ1_comp4CalNComp_calxO),
    .CHQ1_comp3CalPComp_calxO                  (CHQ1_comp3CalPComp_calxO),
    .CHQ1_comp3CalNComp_calxO                  (CHQ1_comp3CalNComp_calxO),
    .CHQ1_comp2CalPComp_calxO                  (CHQ1_comp2CalPComp_calxO),
    .CHQ1_comp2CalNComp_calxO                  (CHQ1_comp2CalNComp_calxO),
    .CHQ1_comp1CalPComp_calxO                  (CHQ1_comp1CalPComp_calxO),
    .CHQ1_comp1CalNComp_calxO                  (CHQ1_comp1CalNComp_calxO),
    .CHQ1_comp0CalPComp_calxO                  (CHQ1_comp0CalPComp_calxO),
    .CHQ1_comp0CalNComp_calxO                  (CHQ1_comp0CalNComp_calxO),
    .CHQ1_compDelayCompDelayxO                 (CHQ1_compDelayCompDelayxO),
    .CHQ1_Fail_detectCH1p1CompFailFlagxI       (CHQ1_Fail_detectCH1p1CompFailFlagxI),
    .CHQ1_Fail_detectCH1p2CompFailFlagxI       (CHQ1_Fail_detectCH1p2CompFailFlagxI),
    .CHQ1_Fail_detectCH1AmpFailFlagxI          (CHQ1_Fail_detectCH1AmpFailFlagxI),
    .CHQ1_SPARESparexO                         (CHQ1_SPARESparexO),
    .CHQ1_N_ValuesNxO                          (CHQ1_N_ValuesNxO),
    .CHQ1_N_ValuesN2xO                         (CHQ1_N_ValuesN2xO),
    .CHQ1_N_ValuesN4xO                         (CHQ1_N_ValuesN4xO),
    .CHQ1_threshold12ThresholdxO               (CHQ1_threshold12ThresholdxO),
    .CHQ1_threshold11ThresholdxO               (CHQ1_threshold11ThresholdxO),
    .CHQ1_threshold10ThresholdxO               (CHQ1_threshold10ThresholdxO),
    .CHQ1_threshold9ThresholdxO                (CHQ1_threshold9ThresholdxO),
    .CHQ1_threshold8ThresholdxO                (CHQ1_threshold8ThresholdxO),
    .CHQ1_threshold7ThresholdxO                (CHQ1_threshold7ThresholdxO),
    .CHQ1_threshold6ThresholdxO                (CHQ1_threshold6ThresholdxO),
    .CHQ1_threshold5ThresholdxO                (CHQ1_threshold5ThresholdxO),
    .CHQ1_threshold4ThresholdxO                (CHQ1_threshold4ThresholdxO),
    .CHQ1_threshold3ThresholdxO                (CHQ1_threshold3ThresholdxO),
    .CHQ1_threshold2ThresholdxO                (CHQ1_threshold2ThresholdxO),
    .CHQ2_calCH2calModexO                      (CHQ2_calCH2calModexO),
    .CHQ2_calShortADCInputxO                   (CHQ2_calShortADCInputxO),
    .CHQ2_calStageCtrlStageDisablexO           (CHQ2_calStageCtrlStageDisablexO),
    .CHQ2_ChannelGainCH2channelGainxO          (CHQ2_ChannelGainCH2channelGainxO),
    .CHQ2_DACN1CH2capControlN1xO               (CHQ2_DACN1CH2capControlN1xO),
    .CHQ2_DACP1CH2capControlP1xO               (CHQ2_DACP1CH2capControlP1xO),
    .CHQ2_DACN2CH2capControlN2xO               (CHQ2_DACN2CH2capControlN2xO),
    .CHQ2_DACP2CH2capControlP2xO               (CHQ2_DACP2CH2capControlP2xO),
    .CHQ2_AMPCH2AmpGainCalPxO                  (CHQ2_AMPCH2AmpGainCalPxO),
    .CHQ2_AMPCH2AmpGainCalNxO                  (CHQ2_AMPCH2AmpGainCalNxO),
    .CHQ2_AMPCH2increaseAmpDelayxO             (CHQ2_AMPCH2increaseAmpDelayxO),
    .CHQ2_MSBCALCH2MSBCalxO                    (CHQ2_MSBCALCH2MSBCalxO),
    .CHQ2_comp12CalPComp_calxO                 (CHQ2_comp12CalPComp_calxO),
    .CHQ2_comp12CalNComp_calxO                 (CHQ2_comp12CalNComp_calxO),
    .CHQ2_comp11CalPComp_calxO                 (CHQ2_comp11CalPComp_calxO),
    .CHQ2_comp11CalNComp_calxO                 (CHQ2_comp11CalNComp_calxO),
    .CHQ2_comp10CalPComp_calxO                 (CHQ2_comp10CalPComp_calxO),
    .CHQ2_comp10CalNComp_calxO                 (CHQ2_comp10CalNComp_calxO),
    .CHQ2_comp9CalPComp_calxO                  (CHQ2_comp9CalPComp_calxO),
    .CHQ2_comp9CalNComp_calxO                  (CHQ2_comp9CalNComp_calxO),
    .CHQ2_comp8CalPComp_calxO                  (CHQ2_comp8CalPComp_calxO),
    .CHQ2_comp8CalNComp_calxO                  (CHQ2_comp8CalNComp_calxO),
    .CHQ2_comp7CalPComp_calxO                  (CHQ2_comp7CalPComp_calxO),
    .CHQ2_comp7CalNComp_calxO                  (CHQ2_comp7CalNComp_calxO),
    .CHQ2_comp6CalPComp_calxO                  (CHQ2_comp6CalPComp_calxO),
    .CHQ2_comp6CalNComp_calxO                  (CHQ2_comp6CalNComp_calxO),
    .CHQ2_comp5CalPComp_calxO                  (CHQ2_comp5CalPComp_calxO),
    .CHQ2_comp5CalNComp_calxO                  (CHQ2_comp5CalNComp_calxO),
    .CHQ2_comp4CalPComp_calxO                  (CHQ2_comp4CalPComp_calxO),
    .CHQ2_comp4CalNComp_calxO                  (CHQ2_comp4CalNComp_calxO),
    .CHQ2_comp3CalPComp_calxO                  (CHQ2_comp3CalPComp_calxO),
    .CHQ2_comp3CalNComp_calxO                  (CHQ2_comp3CalNComp_calxO),
    .CHQ2_comp2CalPComp_calxO                  (CHQ2_comp2CalPComp_calxO),
    .CHQ2_comp2CalNComp_calxO                  (CHQ2_comp2CalNComp_calxO),
    .CHQ2_comp1CalPComp_calxO                  (CHQ2_comp1CalPComp_calxO),
    .CHQ2_comp1CalNComp_calxO                  (CHQ2_comp1CalNComp_calxO),
    .CHQ2_comp0CalPComp_calxO                  (CHQ2_comp0CalPComp_calxO),
    .CHQ2_comp0CalNComp_calxO                  (CHQ2_comp0CalNComp_calxO),
    .CHQ2_compDelayCompDelayxO                 (CHQ2_compDelayCompDelayxO),
    .CHQ2_Fail_detectCH2p1CompFailFlagxI       (CHQ2_Fail_detectCH2p1CompFailFlagxI),
    .CHQ2_Fail_detectCH2p2CompFailFlagxI       (CHQ2_Fail_detectCH2p2CompFailFlagxI),
    .CHQ2_Fail_detectCH2AmpFailFlagxI          (CHQ2_Fail_detectCH2AmpFailFlagxI),
    .CHQ2_SPARESparexO                         (CHQ2_SPARESparexO),
    .CHQ2_N_ValuesNxO                          (CHQ2_N_ValuesNxO),
    .CHQ2_N_ValuesN2xO                         (CHQ2_N_ValuesN2xO),
    .CHQ2_N_ValuesN4xO                         (CHQ2_N_ValuesN4xO),
    .CHQ2_threshold12ThresholdxO               (CHQ2_threshold12ThresholdxO),
    .CHQ2_threshold11ThresholdxO               (CHQ2_threshold11ThresholdxO),
    .CHQ2_threshold10ThresholdxO               (CHQ2_threshold10ThresholdxO),
    .CHQ2_threshold9ThresholdxO                (CHQ2_threshold9ThresholdxO),
    .CHQ2_threshold8ThresholdxO                (CHQ2_threshold8ThresholdxO),
    .CHQ2_threshold7ThresholdxO                (CHQ2_threshold7ThresholdxO),
    .CHQ2_threshold6ThresholdxO                (CHQ2_threshold6ThresholdxO),
    .CHQ2_threshold5ThresholdxO                (CHQ2_threshold5ThresholdxO),
    .CHQ2_threshold4ThresholdxO                (CHQ2_threshold4ThresholdxO),
    .CHQ2_threshold3ThresholdxO                (CHQ2_threshold3ThresholdxO),
    .CHQ2_threshold2ThresholdxO                (CHQ2_threshold2ThresholdxO)
  );

mx_apb_mmap_measADCflags mx_apb_mmap_measADCflags (
    .PClkxCI                                   (PClkxCI),
    .PResetxARBI                               (PResetxARBI),
    .PEnClkxSO                                 (PEnClkxSO_measADCflags),
    .PEnClkxSI                                 (PEnClkxSI),
    .PAddrxDI                                  ({21'h0, PAddrxDI[10:0]}),
    .PSelxSI                                   (PSelxSI_measADCflags),
    .PEnablexSI                                (PEnablexSI),
    .PWritexSI                                 (PWritexSI),
    .PWDataxDI                                 (PWDataxDI),
    .PReadyxSO                                 (PReadyxSO_measADCflags),
    .PRDataxDO                                 (PRDataxDO_measADCflags),
    .PSlverrxSO                                (PSlverrxSO_measADCflags),
    .Adci1Fault_count_ch1stg1_ixI              (Adci1Fault_count_ch1stg1_ixI),
    .Adci1Fault_count_ch1stg2_ixI              (Adci1Fault_count_ch1stg2_ixI),
    .Adci1Fault_count_ch1amp_ixI               (Adci1Fault_count_ch1amp_ixI),
    .Adci2Fault_count_ch2stg1_ixI              (Adci2Fault_count_ch2stg1_ixI),
    .Adci2Fault_count_ch2stg2_ixI              (Adci2Fault_count_ch2stg2_ixI),
    .Adci2Fault_count_ch2amp_ixI               (Adci2Fault_count_ch2amp_ixI),
    .Adcq1Fault_count_ch1stg1_qxI              (Adcq1Fault_count_ch1stg1_qxI),
    .Adcq1Fault_count_ch1stg2_qxI              (Adcq1Fault_count_ch1stg2_qxI),
    .Adcq1Fault_count_ch1amp_qxI               (Adcq1Fault_count_ch1amp_qxI),
    .Adcq2Fault_count_ch2stg1_qxI              (Adcq2Fault_count_ch2stg1_qxI),
    .Adcq2Fault_count_ch2stg2_qxI              (Adcq2Fault_count_ch2stg2_qxI),
    .Adcq2Fault_count_ch2amp_qxI               (Adcq2Fault_count_ch2amp_qxI),
    .Adc_convData_offset_enxO                  (Adc_convData_offset_enxO),
    .Adc_convFault_count_enxO                  (Adc_convFault_count_enxO),
    .Adc_cal_flag_enAdci1EnxO                  (Adc_cal_flag_enAdci1EnxO),
    .Adc_cal_flag_enAdci2EnxO                  (Adc_cal_flag_enAdci2EnxO),
    .Adc_cal_flag_enAdcq1EnxO                  (Adc_cal_flag_enAdcq1EnxO),
    .Adc_cal_flag_enAdcq2EnxO                  (Adc_cal_flag_enAdcq2EnxO)
  );

mx_apb_mmap_measDFE mx_apb_mmap_measDFE (
    .PClkxCI                                   (PClkxCI),
    .PResetxARBI                               (PResetxARBI),
    .PEnClkxSO                                 (PEnClkxSO_measDFE),
    .PEnClkxSI                                 (PEnClkxSI),
    .PAddrxDI                                  ({21'h0, PAddrxDI[10:0]}),
    .PSelxSI                                   (PSelxSI_measDFE),
    .PEnablexSI                                (PEnablexSI),
    .PWritexSI                                 (PWritexSI),
    .PWDataxDI                                 (PWDataxDI),
    .PReadyxSO                                 (PReadyxSO_measDFE),
    .PRDataxDO                                 (PRDataxDO_measDFE),
    .PSlverrxSO                                (PSlverrxSO_measDFE),
    .Padc_gain_ctlPadc_shiftxO                 (Padc_gain_ctlPadc_shiftxO),
    .Padc_gain_ctlPadc_fgain_selxO             (Padc_gain_ctlPadc_fgain_selxO),
    .Padc_gain_ctlPadc_fgain_enxO              (Padc_gain_ctlPadc_fgain_enxO),
    .Padc_gain_ctlMx_swap_iq_enxO              (Padc_gain_ctlMx_swap_iq_enxO),
    .Wb_dcoc_ctlMx_dcoc_est_enxO               (Wb_dcoc_ctlMx_dcoc_est_enxO),
    .Wb_dcoc_ctlMx_dcoc_corr_enxO              (Wb_dcoc_ctlMx_dcoc_corr_enxO),
    .Wb_dcoc_ctlMx_wb_corr_winxO               (Wb_dcoc_ctlMx_wb_corr_winxO),
    .Wb_dcoc_ctlMx_auto_dcoc_enxO              (Wb_dcoc_ctlMx_auto_dcoc_enxO),
    .Wb_dcoc_corr_IMx_dcoc_corr_1_ixO          (Wb_dcoc_corr_IMx_dcoc_corr_1_ixO),
    .Wb_dcoc_corr_IMx_dcoc_corr_2_ixO          (Wb_dcoc_corr_IMx_dcoc_corr_2_ixO),
    .Wb_dcoc_corr_QMx_dcoc_corr_1_qxO          (Wb_dcoc_corr_QMx_dcoc_corr_1_qxO),
    .Wb_dcoc_corr_QMx_dcoc_corr_2_qxO          (Wb_dcoc_corr_QMx_dcoc_corr_2_qxO),
    .Nb_dcoc_ctlMx_dcoc_nb_est_enxO            (Nb_dcoc_ctlMx_dcoc_nb_est_enxO),
    .Nb_dcoc_ctlMx_dcoc_nb_corr_enxO           (Nb_dcoc_ctlMx_dcoc_nb_corr_enxO),
    .Nb_dcoc_ctlMx_nb_corr_winxO               (Nb_dcoc_ctlMx_nb_corr_winxO),
    .Nb_dcoc_ctlMx_auto_dcoc_nb_enxO           (Nb_dcoc_ctlMx_auto_dcoc_nb_enxO),
    .Nb_dcoc_corrMx_dcoc_corr_nb_ixO           (Nb_dcoc_corrMx_dcoc_corr_nb_ixO),
    .Nb_dcoc_corrMx_dcoc_corr_nb_qxO           (Nb_dcoc_corrMx_dcoc_corr_nb_qxO),
    .Adc_imb_ctrlMx_adcimb_corr_enxO           (Adc_imb_ctrlMx_adcimb_corr_enxO),
    .Adc_imb_ctrlMx_adcimb_odden_ixO           (Adc_imb_ctrlMx_adcimb_odden_ixO),
    .Adc_imb_ctrlMx_adcimb_odden_qxO           (Adc_imb_ctrlMx_adcimb_odden_qxO),
    .Adc_imb_ctrlMx_adcimb_corr_ixO            (Adc_imb_ctrlMx_adcimb_corr_ixO),
    .Adc_imb_ctrlMx_adcimb_corr_qxO            (Adc_imb_ctrlMx_adcimb_corr_qxO),
    .Adc_imb_ctrlMx_split_ch_adc_enxO          (Adc_imb_ctrlMx_split_ch_adc_enxO),
    .Wb_iq_corr_ctrlMx_wb_corr_est_enxO        (Wb_iq_corr_ctrlMx_wb_corr_est_enxO),
    .Wb_iq_corr_ctrlMx_iqcorr_enxO             (Wb_iq_corr_ctrlMx_iqcorr_enxO),
    .Wb_iq_corr_ctrlMx_iqcorr_1xO              (Wb_iq_corr_ctrlMx_iqcorr_1xO),
    .Wb_iq_corr_ctrlMx_iqcorr_2xO              (Wb_iq_corr_ctrlMx_iqcorr_2xO),
    .Nb_iq_corr_ctrlMx_nb_corr_est_enxO        (Nb_iq_corr_ctrlMx_nb_corr_est_enxO),
    .Nb_iq_corr_ctrlMx_iqcorr_nb_enxO          (Nb_iq_corr_ctrlMx_iqcorr_nb_enxO),
    .Nb_iq_corr_ctrlMx_iqcorr_nb_1xO           (Nb_iq_corr_ctrlMx_iqcorr_nb_1xO),
    .Nb_iq_corr_ctrlMx_iqcorr_nb_2xO           (Nb_iq_corr_ctrlMx_iqcorr_nb_2xO),
    .Init_sample_ctrlMx_data_w_chopxO          (Init_sample_ctrlMx_data_w_chopxO),
    .Hist_ctrlHist_count_enxO                  (Hist_ctrlHist_count_enxO),
    .Hist_ctrlHist_absbin_enxO                 (Hist_ctrlHist_absbin_enxO),
    .Hist_ctrlHist_count_clrxO                 (Hist_ctrlHist_count_clrxO),
    .Hist_ctrlHist_max_countxO                 (Hist_ctrlHist_max_countxO),
    .Filts_ctrl_1Filts_enxO                    (Filts_ctrl_1Filts_enxO),
    .Filts_ctrl_1Init_ds_ratexO                (Filts_ctrl_1Init_ds_ratexO),
    .Filts_ctrl_2Fr_offset_ixO                 (Filts_ctrl_2Fr_offset_ixO),
    .Filts_ctrl_2Fr_offset_qxO                 (Filts_ctrl_2Fr_offset_qxO),
    .Filts_ctrl_2Mx_farrow_gain_selxO          (Filts_ctrl_2Mx_farrow_gain_selxO),
    .Filts_ctrl_3Fr_ctrlxO                     (Filts_ctrl_3Fr_ctrlxO),
    .Wb_dcoc_est_iDcoc_estimate_1_ixI          (Wb_dcoc_est_iDcoc_estimate_1_ixI),
    .Wb_dcoc_est_iDcoc_estimate_2_ixI          (Wb_dcoc_est_iDcoc_estimate_2_ixI),
    .Wb_dcoc_est_qDcoc_estimate_1_qxI          (Wb_dcoc_est_qDcoc_estimate_1_qxI),
    .Wb_dcoc_est_qDcoc_estimate_2_qxI          (Wb_dcoc_est_qDcoc_estimate_2_qxI),
    .Nb_dcoc_estsDcoc_estimate_nb_ixI          (Nb_dcoc_estsDcoc_estimate_nb_ixI),
    .Nb_dcoc_estsDcoc_estimate_nb_qxI          (Nb_dcoc_estsDcoc_estimate_nb_qxI),
    .Mx_statusDcoc_count_donexI                (Mx_statusDcoc_count_donexI),
    .Mx_statusCorr_count_donexI                (Mx_statusCorr_count_donexI),
    .Mx_statusHist_overflowxI                  (Mx_statusHist_overflowxI),
    .Mx_statusHist_count_donexI                (Mx_statusHist_count_donexI),
    .Mx_statusDcoc_count_nb_donexI             (Mx_statusDcoc_count_nb_donexI),
    .Mx_statusCorr_count_nb_donexI             (Mx_statusCorr_count_nb_donexI),
    .Wb_pwrMx_wb_pwrxI                         (Wb_pwrMx_wb_pwrxI),
    .Nb_pwrMx_nb_pwrxI                         (Nb_pwrMx_nb_pwrxI),
    .Corr_iwbCorr_iwb_outxI                    (Corr_iwbCorr_iwb_outxI),
    .Corr_qwbCorr_qwb_outxI                    (Corr_qwbCorr_qwb_outxI),
    .Corr_iqwbCorr_iqwb_outxI                  (Corr_iqwbCorr_iqwb_outxI),
    .Corr_inbCorr_inb_outxI                    (Corr_inbCorr_inb_outxI),
    .Corr_qnbCorr_qnb_outxI                    (Corr_qnbCorr_qnb_outxI),
    .Corr_iqnbCorr_iqnb_outxI                  (Corr_iqnbCorr_iqnb_outxI),
    .Corr_iwb_1Corr_iwb_1_outxI                (Corr_iwb_1Corr_iwb_1_outxI),
    .Corr_iwb_2Corr_iwb_2_outxI                (Corr_iwb_2Corr_iwb_2_outxI),
    .Corr_qwb_1Corr_qwb_1_outxI                (Corr_qwb_1Corr_qwb_1_outxI),
    .Corr_qwb_2Corr_qwb_2_outxI                (Corr_qwb_2Corr_qwb_2_outxI),
    .Hist_i_0Hist_out_i_0xI                    (Hist_i_0Hist_out_i_0xI),
    .Hist_i_0Hist_out_i_1xI                    (Hist_i_0Hist_out_i_1xI),
    .Hist_i_1Hist_out_i_2xI                    (Hist_i_1Hist_out_i_2xI),
    .Hist_i_1Hist_out_i_3xI                    (Hist_i_1Hist_out_i_3xI),
    .Hist_i_2Hist_out_i_4xI                    (Hist_i_2Hist_out_i_4xI),
    .Hist_i_2Hist_out_i_5xI                    (Hist_i_2Hist_out_i_5xI),
    .Hist_i_3Hist_out_i_6xI                    (Hist_i_3Hist_out_i_6xI),
    .Hist_i_3Hist_out_i_7xI                    (Hist_i_3Hist_out_i_7xI),
    .Hist_i_4Hist_out_i_8xI                    (Hist_i_4Hist_out_i_8xI),
    .Hist_i_4Hist_out_i_9xI                    (Hist_i_4Hist_out_i_9xI),
    .Hist_i_5Hist_out_i_10xI                   (Hist_i_5Hist_out_i_10xI),
    .Hist_i_5Hist_out_i_11xI                   (Hist_i_5Hist_out_i_11xI),
    .Hist_i_6Hist_out_i_12xI                   (Hist_i_6Hist_out_i_12xI),
    .Hist_i_6Hist_out_i_13xI                   (Hist_i_6Hist_out_i_13xI),
    .Hist_i_7Hist_out_i_14xI                   (Hist_i_7Hist_out_i_14xI),
    .Hist_i_7Hist_out_i_15xI                   (Hist_i_7Hist_out_i_15xI),
    .Hist_i_8Hist_out_i_16xI                   (Hist_i_8Hist_out_i_16xI),
    .Hist_i_8Hist_out_i_17xI                   (Hist_i_8Hist_out_i_17xI),
    .Hist_i_9Hist_out_i_18xI                   (Hist_i_9Hist_out_i_18xI),
    .Hist_i_9Hist_out_i_19xI                   (Hist_i_9Hist_out_i_19xI),
    .Hist_i_10Hist_out_i_20xI                  (Hist_i_10Hist_out_i_20xI),
    .Hist_i_10Hist_out_i_21xI                  (Hist_i_10Hist_out_i_21xI),
    .Hist_i_11Hist_out_i_22xI                  (Hist_i_11Hist_out_i_22xI),
    .Hist_i_11Hist_out_i_23xI                  (Hist_i_11Hist_out_i_23xI),
    .Hist_i_12Hist_out_i_24xI                  (Hist_i_12Hist_out_i_24xI),
    .Hist_i_12Hist_out_i_25xI                  (Hist_i_12Hist_out_i_25xI),
    .Hist_i_13Hist_out_i_26xI                  (Hist_i_13Hist_out_i_26xI),
    .Hist_i_13Hist_out_i_27xI                  (Hist_i_13Hist_out_i_27xI),
    .Hist_i_14Hist_out_i_28xI                  (Hist_i_14Hist_out_i_28xI),
    .Hist_i_14Hist_out_i_29xI                  (Hist_i_14Hist_out_i_29xI),
    .Hist_i_15Hist_out_i_30xI                  (Hist_i_15Hist_out_i_30xI),
    .Hist_i_15Hist_out_i_31xI                  (Hist_i_15Hist_out_i_31xI),
    .Hist_q_0Hist_out_i_0xI                    (Hist_q_0Hist_out_i_0xI),
    .Hist_q_0Hist_out_i_1xI                    (Hist_q_0Hist_out_i_1xI),
    .Hist_q_1Hist_out_i_2xI                    (Hist_q_1Hist_out_i_2xI),
    .Hist_q_1Hist_out_i_3xI                    (Hist_q_1Hist_out_i_3xI),
    .Hist_q_2Hist_out_i_4xI                    (Hist_q_2Hist_out_i_4xI),
    .Hist_q_2Hist_out_i_5xI                    (Hist_q_2Hist_out_i_5xI),
    .Hist_q_3Hist_out_i_6xI                    (Hist_q_3Hist_out_i_6xI),
    .Hist_q_3Hist_out_i_7xI                    (Hist_q_3Hist_out_i_7xI),
    .Hist_q_4Hist_out_i_8xI                    (Hist_q_4Hist_out_i_8xI),
    .Hist_q_4Hist_out_i_9xI                    (Hist_q_4Hist_out_i_9xI),
    .Hist_q_5Hist_out_i_10xI                   (Hist_q_5Hist_out_i_10xI),
    .Hist_q_5Hist_out_i_11xI                   (Hist_q_5Hist_out_i_11xI),
    .Hist_q_6Hist_out_i_12xI                   (Hist_q_6Hist_out_i_12xI),
    .Hist_q_6Hist_out_i_13xI                   (Hist_q_6Hist_out_i_13xI),
    .Hist_q_7Hist_out_i_14xI                   (Hist_q_7Hist_out_i_14xI),
    .Hist_q_7Hist_out_i_15xI                   (Hist_q_7Hist_out_i_15xI),
    .Hist_q_8Hist_out_i_16xI                   (Hist_q_8Hist_out_i_16xI),
    .Hist_q_8Hist_out_i_17xI                   (Hist_q_8Hist_out_i_17xI),
    .Hist_q_9Hist_out_i_18xI                   (Hist_q_9Hist_out_i_18xI),
    .Hist_q_9Hist_out_i_19xI                   (Hist_q_9Hist_out_i_19xI),
    .Hist_q_10Hist_out_i_20xI                  (Hist_q_10Hist_out_i_20xI),
    .Hist_q_10Hist_out_i_21xI                  (Hist_q_10Hist_out_i_21xI),
    .Hist_q_11Hist_out_i_22xI                  (Hist_q_11Hist_out_i_22xI),
    .Hist_q_11Hist_out_i_23xI                  (Hist_q_11Hist_out_i_23xI),
    .Hist_q_12Hist_out_i_24xI                  (Hist_q_12Hist_out_i_24xI),
    .Hist_q_12Hist_out_i_25xI                  (Hist_q_12Hist_out_i_25xI),
    .Hist_q_13Hist_out_i_26xI                  (Hist_q_13Hist_out_i_26xI),
    .Hist_q_13Hist_out_i_27xI                  (Hist_q_13Hist_out_i_27xI),
    .Hist_q_14Hist_out_i_28xI                  (Hist_q_14Hist_out_i_28xI),
    .Hist_q_14Hist_out_i_29xI                  (Hist_q_14Hist_out_i_29xI),
    .Hist_q_15Hist_out_i_30xI                  (Hist_q_15Hist_out_i_30xI),
    .Hist_q_15Hist_out_i_31xI                  (Hist_q_15Hist_out_i_31xI),
    .Adc_tmodeTmodexO                          (Adc_tmodeTmodexO)
  );
endmodule
